module ternary_min(a[1:0], b[1:0], out[1:0]);
  input [1:0] a
  input [1:0] b;
  output [1:0] out;
  // TODO: implementation
endmodule

module ternary_max(a[1:0], b[1:0], out[1:0]);
  input [1:0] a
  input [1:0] b;
  output [1:0] out;
  // TODO: implementation
endmodule

module ternary_any(a[1:0], b[1:0], out[1:0]);
  input [1:0] a
  input [1:0] b;
  output [1:0] out;
  // TODO: implementation
endmodule

module ternary_consensus(a[1:0], b[1:0], out[1:0]);
  input [1:0] a
  input [1:0] b;
  output [1:0] out;
  // TODO: implementation
endmodule
